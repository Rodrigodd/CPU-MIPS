module MUX(
	input clk, rst
);
endmodule

