module ALU(
	input clk, rst
);
endmodule

