module ADDRDecoding(
	input clk, rst,
	input [31:0] addr,
	output cs
);

endmodule

