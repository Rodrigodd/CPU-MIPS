module Extend(
	input clk, rst,
	input [31:0] instr,
	output [31:0] imm
);

endmodule

