module Control(
	input clk, rst
);
endmodule

