module InstructionMemory(
	input clk, rst,
	input [31:0] addr,
	output [31:0] data
);
endmodule

