module DataMemory(
	input clk, rst
);
endmodule

