module Extend(
	input clk, rst
);
endmodule

