module Control(
	input clk, rst,
	input [31:0] instr,
	output [4:0] a_reg, b_reg,
	output [10:0] ctrl_ex
);
endmodule

