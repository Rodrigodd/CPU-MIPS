module Register(
	input clk, rst
);
endmodule

