module InstructionMemory(
	input clk, rst
);
endmodule

