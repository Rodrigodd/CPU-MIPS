module ADDRDecoding(
	input clk, rst
);
endmodule

