module Multiplicador(
	input clk, rst
);
endmodule

