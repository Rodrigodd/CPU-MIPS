module ALU(
	input clk, rst,
	input [31:0] a, c_ex,
	input [1:0] op_sel,
	output [31:0] op
);
endmodule

