module PLL(
	input clk, rst
);
endmodule

