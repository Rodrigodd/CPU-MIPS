module PC(
	input clk, rst
);
endmodule

