module RegisterFile(
	input clk, rst
);
endmodule

